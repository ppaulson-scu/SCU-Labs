*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'ppaulson' on Tue May 16 2017 at 15:23:31

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $UpdatedFiles/default.group/logic.views/153OR
*
.subckt 153OR  OUT A B

        M3 N$12 A GROUND GROUND N L=.4u W=1.2u M=1
        M1 N$12 B GROUND GROUND N L=.4u W=1.2u M=1
        M6 OUT N$12 VDD VDD P L=.4u W=2.4u M=1
        M5 OUT N$12 GROUND GROUND N L=.4u W=1.2u M=1
        M4 N$12 B N$8 VDD P L=.4u W=4.8u M=1
        M2 N$8 A VDD VDD P L=.4u W=4.8u M=1
.ends 153OR

*
* Component pathname : $UpdatedFiles/default.group/logic.views/inverter
*
.subckt INVERTER  OUT IN

        M2 OUT IN VDD VDD P L=0.4u W=3.6u M=1
        M1 OUT IN GROUND GROUND N L=0.4u W=1.2u M=1
.ends INVERTER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/153XOR
*
.subckt 153XOR  XOR A B

        X_INVERTER1 XOR N$3 INVERTER
        M2 B A N$3 GROUND N L=0.4u W=1.2u M=2
        M4 A B N$3 GROUND N L=0.4u W=1.2u M=2
        M3 N$3 B N$2 VDD P L=0.4u W=2.4u M=2
        M1 N$2 A VDD VDD P L=0.4u W=2.4u M=2
.ends 153XOR

*
* Component pathname : $UpdatedFiles/default.group/logic.views/153AND
*
.subckt 153AND  OUT A B

        M1 OUT N$4 GROUND GROUND N L=.4u W=1.2u M=1
        M3 N$6 A GROUND GROUND N L=.4u W=2.4u M=1
        M5 N$4 B N$6 GROUND N L=.4u W=2.4u M=1
        M4 N$4 B VDD VDD P L=.4u W=2.4u M=1
        M6 N$4 A VDD VDD P L=.4u W=2.4u M=1
        M2 OUT N$4 VDD VDD P L=.4u W=2.4u M=1
.ends 153AND

*
* Component pathname : $UpdatedFiles/default.group/logic.views/HalfAdder
*
.subckt HALFADDER  C S X Y

        X_153XOR1 S Y X 153XOR
        X_153AND1 C X Y 153AND
.ends HALFADDER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/FullAdder
*
.subckt FULLADDER  C+1 S A B C

        X_153OR1 C+1 N$205 N$203 153OR
        X_HALFADDER2 N$205 S N$204 C HALFADDER
        X_HALFADDER1 N$203 N$204 A B HALFADDER
.ends FULLADDER

*
* Component pathname : $UpdatedFiles/default.group/logic.views/4BitAdder
*
.subckt 4BITADDER  COUT S0 S1 S2 S3 A0 A1 A2 A3 B0 B1 B2 B3 CIN

        X_FULLADDER4 COUT S3 B3 A3 N$6 FULLADDER
        X_FULLADDER3 N$6 S2 B2 A2 N$4 FULLADDER
        X_FULLADDER2 N$4 S1 B1 A1 N$2 FULLADDER
        X_FULLADDER1 N$2 S0 A0 B0 CIN FULLADDER
.ends 4BITADDER

*
* MAIN CELL: Component pathname : $UpdatedFiles/default.group/logic.views/Test
*
        V9 VDD GROUND DC 5V
        V7 N$5 GROUND PATTERN 5 0 0 1n 1n 50n 11010010110
        V8 N$1 GROUND PATTERN 5 0 0 1n 1n 50n 00110011001
        V6 N$6 GROUND PATTERN 5 0 0 1n 1n 50n 01010111101
        V5 N$7 GROUND PATTERN 5 0 0 1n 1n 50n 11111101010
        V3 N$2 GROUND PATTERN 5 0 0 1n 1n 50n 01011010010
        V4 N$4 GROUND PATTERN 5 0 0 1n 1n 50n 01100110011
        V2 N$3 GROUND PATTERN 5 0 0 1n 1n 50n 01010000101
        V1 N$13 GROUND PATTERN 5 0 0 1n 1n 50n 00000101010
        X_4BITADDER1 COUT S0 S1 S2 S3 N$1 N$2 N$3 N$13 N$4 N$5 N$6 N$7 GROUND 4BITADDER
*
.end
